* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
R1 1 0 21.58680303547402
C2 1 2 2.1373072312350514
R2 2 0 0.2158464457101714
C3 2 3 0.021586781448670544
R3 3 0 0.00215868028218085
C4 3 4 0.0002158680281306431
R4 4 0 2.1586825060555236e-05
C5 4 5 2.1584600529665642e-06
R5 5 0 2.180707631106713e-07
R6 5 0 2.180707631106713e-07
.AC DEC 100 1 1000000
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
