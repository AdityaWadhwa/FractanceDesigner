* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
R1 1 2 5.372181010131195
C1 1 2 1.0124379632299796
R2 2 3 0.06569539305200849
C2 2 3 2.3413349529430585
R3 3 4 0.002654093879301143
C3 3 4 1.6389344670601411
R4 4 5 0.00010722539272376618
C4 4 5 1.1472541269420988
R5 5 6 4.3319058660401535e-06
C5 5 6 0.8030778888594693
R6 6 7 1.7500899698802218e-07
C6 6 7 0.5621545222016285
R7 7 8 7.070363478316096e-09
C7 7 8 0.39350816554114004
R8 8 9 2.856426845239703e-10
C8 8 9 0.2754557158787981
R9 9 10 1.1539964454768398e-11
C9 9 10 0.19281900111515865
R10 10 11 2.331072819863216e-13
C10 10 11 0.26994660156122213
R11 11 0 1.4528681480519884e-13
.AC DEC 100 1.0 1000000.0
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
