* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
R1 1 2 1.5310955542480119e-06
C1 1 2 0.08170613604718352
R2 2 3 1.6132026470174018e-05
C2 2 3 0.13790119903731643
R3 3 4 0.0001617808927558726
C3 3 4 0.24452864461254412
R4 4 5 0.0016180760852820904
C4 4 5 0.4347684581624912
R5 5 6 0.01618236290835089
C5 5 6 0.7730632563682562
R6 6 7 0.16208316335844217
C6 6 7 1.3725212088926397
R7 7 8 1.6684677425936003
C7 7 8 2.3710414903380594
R8 8 9 35.97878894226995
C8 8 9 1.9552866160016769
R9 9 0 3.7827320109503437e-07
.AC DEC 100 1 1000
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
