* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
R1 1 2 0.037037037037037035
C2 2 0 0.11126373626373627
R2 2 3 0.18595146871008938
C3 3 0 0.2614182692307693
R3 3 4 0.33799874256420204
C4 4 0 0.41605184366414827
R4 4 5 0.49596993617886226
C5 5 0 0.5781896945038527
R5 5 6 0.6632056058100293
C6 6 0 0.7515871183185393
R6 6 7 0.844000924330203
C7 7 0 0.9412405506158444
R7 7 8 1.04426650792174
C8 8 0 1.154261995106964
R8 8 9 1.2727120516811063
C9 9 0 1.4015190288911366
R9 9 10 1.5431761204022223
C10 10 0 1.7010372084528238
R10 10 11 1.879753628144543
C11 11 0 2.086015738160563
R11 11 12 2.329887681051604
C12 12 0 2.6273917955626938
R12 12 13 3.0060074013371145
C13 13 0 3.51795540998879
R13 13 0 9.081329549427794
.AC DEC 1 0.1 100
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
