* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
R1 1 2 0.0006453982796935868
C1 1 2 0.014406180581533857
R2 2 3 0.0012725681893588031
C2 2 3 0.018352515305238
R3 3 4 0.002157068594297493
C3 3 4 0.027196480278422495
R4 4 5 0.003503689681596965
C4 4 5 0.04205823309850728
R5 5 6 0.005605777249781898
C5 5 6 0.06602992760319268
R6 6 7 0.00891768241704329
C6 6 7 0.10426166496473913
R7 7 8 0.014154442786600132
C7 7 8 0.1649999757975353
R8 8 9 0.022446504754539368
C8 8 9 0.26135326691410093
R9 9 10 0.035583931393574963
C9 9 10 0.4141166857129336
R10 10 11 0.0564032732824955
C10 10 11 0.6562545831495191
R11 11 12 0.08940169274404411
C11 11 12 1.0399941968544693
R12 12 13 0.1417150418238487
C12 12 13 1.6480132857877168
R13 13 14 0.2246874903852943
C13 13 14 2.610945245924333
R14 14 15 0.35643744274422945
C14 14 15 4.134217668012565
R15 15 16 0.5662395600004663
C15 15 16 6.536969369685508
R16 16 17 0.9027630903485048
C16 16 17 10.299185094826791
R17 17 18 1.4526756963913008
C17 17 18 16.077110142466207
R18 18 19 2.396742642878488
C18 18 19 24.476834698263556
R19 19 20 4.268827671384615
C19 19 20 34.519781232031484
R20 20 21 11.034463689840457
C20 20 21 33.54481707194572
R21 21 0 0.002158680303547402
.AC DEC 100 1 1000
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
