* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
R1 1 2 38.86550831153718
C1 1 2 45.696044568978316
R2 2 3 9.769150837043831
C2 2 3 29.087482089281323
R3 3 4 3.9076603348175327
C3 3 4 11.63499283571253
R4 4 5 1.5630641339270133
C4 4 5 4.653997134285012
R5 5 6 0.6252256535708053
C5 5 6 1.861598853714005
R6 6 7 0.25009026142832214
C6 6 7 0.744639541485602
R7 7 8 0.10003610457132886
C7 7 8 0.2978558165942408
R8 8 9 0.04001444182853154
C8 8 9 0.11914232663769633
R9 9 10 0.01600577673141262
C9 9 10 0.04765693065507854
R10 10 11 0.0064023106925650474
C10 10 11 0.019062772262031416
R11 11 12 0.0025609242770260193
C11 11 12 0.007625108904812567
R12 12 13 0.0005121848554052039
C12 12 13 0.006100087123850053
R13 13 0 0.0011179527143259334
.AC DEC 100 0.001 1000.0
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
