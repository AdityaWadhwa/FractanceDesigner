* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
R1 1 2 2.3291
C1 1 2 1.1914
R2 2 3 0.23786
C2 2 3 1.1573
R3 3 4 0.047192
C3 3 4 0.57865
R4 4 5 0.0093629
C4 4 5 0.28933
R5 5 6 0.0018576
C5 5 6 0.14466
R6 6 7 0.00036855
C6 6 7 0.072331
R7 7 8 7.312e-05
C7 7 8 0.036166
R8 8 9 1.4507e-05
C8 8 9 0.018083
R9 9 10 2.8782e-06
C9 9 10 0.0090414
R10 10 11 5.7103e-07
C10 10 11 0.0045207
R11 11 12 1.1329e-07
C11 11 12 0.0022604
R12 12 13 1.1239e-08
C12 12 13 0.0022604
R13 13 0 1.3897e-08
.AC DEC 100 1 1000000
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
