['* Matlab created *.cir-file *']
['.lib C:\\Cadence\\SPB_17.2\\tools\\pspice\\library\\eval.lib']
['VIN        1   0   AC 1V']
['R1 1 2 0.004466465413723158']
['C1 2 0 0.1699293784879202']
['R2 1 3 0.10944709326979155']
['C2 3 0 0.10067326662828437']
['R3 1 4 0.3943572830972851']
['C3 4 0 0.09077568318875885']
['R4 1 5 0.8799657438081956']
['C4 5 0 0.09536431612559092']
['R5 1 6 1.5634964067290835']
['C5 6 0 0.11375807385553609']
['R6 1 7 2.4395272615944728']
['C6 7 0 0.15705717488835863']
['R7 1 8 3.550428299268764']
['C7 8 0 0.2695097724763911']
['R8 1 9 5.208383208325146']
['C8 9 0 0.7330618273265841']
['R9 1 9 18.181590757812568']
['.AC DEC 100 0.01 100']
['.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)']
['.END']
