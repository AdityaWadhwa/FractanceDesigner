* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
R1 1 0 56.2341
C2 1 2 1.1197
R2 2 0 6.3569
C3 2 3 0.99302
R3 3 0 1.3405
C4 3 4 0.52082
R4 4 0 0.2723
C5 4 5 0.25453
R5 5 0 0.060977
C6 5 6 0.095029



R7 6 0 0.028376
.AC DEC 100 0.01 1000
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
