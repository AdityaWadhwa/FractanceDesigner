* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
Rp 1 0 21.24298386366024
Cp 1 0 0.002414529118663077
R1 1 2 3.681605899141823
C1 2 0 4.322976099342793
R2 1 3 0.5438092311884086
C2 3 0 0.6385458882433493
R3 1 4 0.08032594689036705
C3 4 0 0.09431947853111548
.AC DEC 100 0.01 100
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
