* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
Rp 1 0 0.9957082169652448
Cp 1 0 7.977991014899577e-05
R1 1 2 0.7501342587565025
C1 2 0 0.2121686101308404
R2 1 3 0.32230938013324567
C2 3 0 0.09116225851138098
R3 1 4 0.13848632469350816
C3 4 0 0.03916958956261668
R4 1 5 0.05950327017844535
C4 5 0 0.016829955417485713
R5 1 6 0.025566706097263043
C5 6 0 0.007231308842329232
R6 1 7 0.010985219109866835
C6 7 0 0.0031070686924589003
R7 1 8 0.004720007279494716
C7 8 0 0.0013350108631992423
R8 1 9 0.0020280404510523388
C8 9 0 0.0005736126816847199
R9 1 10 0.0008713859592913322
C9 10 0 0.00024646354397524467
.AC DEC 100 1.0 1000000.0
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
