* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
Rp 1 0 31.48705850555284
Cp 1 0 0.0025228622759440986
R1 1 2 23.721328085926544
C1 2 0 6.70936056005731
R2 1 3 10.19231752458081
C2 3 0 2.8828037354103473
R3 1 4 4.3793221081710545
C3 4 0 1.2386511803182723
R4 1 5 1.8816586199226109
C4 5 0 0.5322099203834486
R5 1 6 0.8084902353546563
C5 6 0 0.22867406405875793
R6 1 7 0.34738312983186664
C6 7 0 0.09825413914771355
R7 1 8 0.14925973575778267
C7 8 0 0.04221675028777068
R8 1 9 0.06413227012280615
C8 9 0 0.018139225688808654
R9 1 10 0.02755564352451373
C9 10 0 0.00779386159158843
.AC DEC 100 0.001 1000.0
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
