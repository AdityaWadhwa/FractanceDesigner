* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
R1 1 2 0.02202
C1 2 0 0.020436
R2 1 3 0.11891
C2 3 0 0.01041
R3 1 4 0.16627
C3 4 0 0.026647
R4 1 5 0.31086
C4 5 0 0.051011
R5 1 6 0.58721
C5 6 0 0.096653
R6 1 7 1.1106
C6 7 0 0.18291
R7 1 8 2.1008
C7 8 0 0.34608
R8 1 9 3.9742
C8 9 0 0.65476
R9 1 10 7.5174
C9 10 0 1.2389
R10 1 11 14.2153
C10 11 0 2.3449
R11 1 12 26.8683
C11 12 0 4.4403
R12 1 13 51.325
C12 13 0 8.3195
R13 1 14 45.4125
C13 14 0 48.9341

R14 1 14 0.015
.AC DEC 100 0.001 1000
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
