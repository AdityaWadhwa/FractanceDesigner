* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
R1 1 0 682.6346
C2 1 2 308.0689































R3 2 0 234.5829
.AC DEC 100 0.001 1000
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
