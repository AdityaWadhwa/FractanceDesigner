* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
R1 1 2 0.037037
C2 2 0 0.11126
R2 2 3 0.18595
C3 3 0 0.26142
R3 3 4 0.338
C4 4 0 0.41605
R4 4 5 0.49597
C5 5 0 0.57819
R5 5 6 0.66321
C6 6 0 0.75159
R6 6 7 0.844
C7 7 0 0.94124
R7 7 8 1.0443
C8 8 0 1.1543
R8 8 9 1.2727
C9 9 0 1.4015
R9 9 10 1.5432
C10 10 0 1.701
R10 10 11 1.8798
C11 11 0 2.086
R11 11 12 2.3299
C12 12 0 2.6274
R12 12 13 3.006
C13 13 0 3.518
R13 13 14 4.2787
C14 14 0 5.6159



R15 14 0 9.0813
.AC DEC 100 0.1 10
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
