* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
R1 1 2 1.5198898948036383
C1 1 2 1.1685056964139169
R2 2 3 0.24163793769988043
C2 2 3 0.743803732604398
R3 3 4 0.061134398238069744
C3 3 4 0.29752149304175923
R4 4 5 0.015467002754231645
C4 4 5 0.1190085972167037
R5 5 6 0.0039131516968206066
C5 5 6 0.047603438886681476
R6 6 7 0.0009900273792956135
C6 6 7 0.019041375554672592
R7 7 8 0.00025047692696179017
C7 7 8 0.0076165502218690385
R8 8 9 6.337066252133292e-05
C8 8 9 0.003046620088747615
R9 9 10 1.603277761789723e-05
C9 9 10 0.0012186480354990463
R10 10 11 4.056292737327999e-06
C10 10 11 0.0004874592141996185
R11 11 12 1.0262420625439837e-06
C11 11 12 0.0001949836856798474
R12 12 13 1.2981962091181395e-07
C12 12 13 0.00015598694854387793
R13 13 0 1.8891567562630236e-07
.AC DEC 100 1 1000000
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
