['* Matlab created *.cir-file *']
['.lib C:\\Cadence\\SPB_17.2\\tools\\pspice\\library\\eval.lib']
['VIN        1   0   AC 1V']
['R1 1 2 0.06838811614413393']
['C1 2 0 0.06580223849427881']
['R2 1 3 0.5930756494431398']
['C2 3 0 0.018798421933769564']
['R3 1 4 0.6125322543737914']
['C3 4 0 0.04286061823867516']
['R4 1 5 0.916851535021896']
['C4 5 0 0.0674286220402618']
['R5 1 6 1.401323840869538']
['C5 6 0 0.10388687861148668']
['R6 1 7 2.1484239204240163']
['C6 7 0 0.15956408150578677']
['R7 1 8 3.2958596666895392']
['C7 8 0 0.2449301855020474']
['R8 1 9 5.056752354163437']
['C8 9 0 0.3759198383044014']
['R9 1 10 7.758618000705936']
['C9 10 0 0.5769503859509636']
['R10 1 11 11.908508249408259']
['C10 11 0 0.8851591914896837']
['R11 1 12 18.34712887852123']
['C11 12 0 1.3529026298978373']
['R12 1 13 29.36346517590909']
['C12 13 0 1.990596585431996']
['R13 1 14 14.622423549327197']
['C13 14 0 15.197051390384479']
['R14 1 14 0.04743416490252569']
['.AC DEC 100 0.01 100']
['.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)']
['.END']
