* Matlab created *.cir-file *
.lib C:\Cadence\SPB_17.2\tools\pspice\library\eval.lib
VIN        1   0   AC 1V
R1 1 2 60.4142
C1 1 2 4.5933
R2 2 3 6.1699
C2 2 3 4.4617
R3 3 4 1.2241
C3 3 4 2.2308
R4 4 5 0.24286
C4 4 5 1.1154
R5 5 6 0.048184
C5 5 6 0.55771
R6 6 7 0.0095597
C6 6 7 0.27886
R7 7 8 0.0018966
C7 7 8 0.13943
R8 8 9 0.00037629
C8 8 9 0.069714
R9 9 10 7.4656e-05
C9 9 10 0.034857
R10 10 11 1.4812e-05
C10 10 11 0.017428
R11 11 12 2.9387e-06
C11 11 12 0.0087142
R12 12 13 2.9152e-07
C12 12 13 0.0087142
R13 13 0 3.6046e-07
.AC DEC 100 0.01 1000
.PRINT AC VM(1) VP(1) IM(VIN) IP(VIN)
.END
